(* vim:ft=coq *)

(* `Require Export` statement to tell Rocq to use the String module from the standard library *)
From Stdlib Require Export String.
